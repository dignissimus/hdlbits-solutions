module top_module(output onex);
    assign one = 1;
endmodule

