module top_module(input a, input b, output out);
	mod_a module_instance(.in1(a), .in2(b), .out(out));
endmodule
